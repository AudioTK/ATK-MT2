*
Vin	Vin	0	AC	1
Vdd Vdd	0	DC -4.5
Vcc	Vcc	0	DC 4.5
*
*	V-	V+	Vout
Z1	2	Vin	Vout
R030	2	Vout	3.3k
C022	2	Vout	47p

* Gyrator
C020	2	3	0.022u
R027	3	4	470
R024	4	Vdd	10k
C017	3	5	0.047u
R025	0	5	470k
Q007	Vcc	5	4	trans

* Gyrator
C024	2	6	0.015u
R034	6	7	1k
R037	7	Vdd	10k
C025	6	8	0.0015u
R036	0	8	47k
Q008	Vcc	8	7	trans

.model trans npn(vt=26e-3 is=1e-12 ne=1 br=1 bf=100)
